module PDPW16KD_wrapper2 (
	input wire JADA0_EBR,
	input wire JADA10_EBR,
	input wire JADA11_EBR,
	input wire JADA12_EBR,
	input wire JADA13_EBR,
	input wire JADA1_EBR,
	input wire JADA2_EBR,
	input wire JADA3_EBR,
	input wire JADA4_EBR,
	input wire JADA5_EBR,
	input wire JADA6_EBR,
	input wire JADA7_EBR,
	input wire JADA8_EBR,
	input wire JADA9_EBR,
	input wire JADB0_EBR,
	input wire JADB10_EBR,
	input wire JADB11_EBR,
	input wire JADB12_EBR,
	input wire JADB13_EBR,
	input wire JADB1_EBR,
	input wire JADB2_EBR,
	input wire JADB3_EBR,
	input wire JADB4_EBR,
	input wire JADB5_EBR,
	input wire JADB6_EBR,
	input wire JADB7_EBR,
	input wire JADB8_EBR,
	input wire JADB9_EBR,
	input wire JCEA_EBR,
	input wire JCEB_EBR,
	input wire JCLKA_EBR,
	input wire JCLKB_EBR,
	input wire JCSA0_EBR,
	input wire JCSA1_EBR,
	input wire JCSA2_EBR,
	input wire JCSB0_EBR,
	input wire JCSB1_EBR,
	input wire JCSB2_EBR,
	input wire JDIA0_EBR,
	input wire JDIA10_EBR,
	input wire JDIA11_EBR,
	input wire JDIA12_EBR,
	input wire JDIA13_EBR,
	input wire JDIA14_EBR,
	input wire JDIA15_EBR,
	input wire JDIA16_EBR,
	input wire JDIA17_EBR,
	input wire JDIA1_EBR,
	input wire JDIA2_EBR,
	input wire JDIA3_EBR,
	input wire JDIA4_EBR,
	input wire JDIA5_EBR,
	input wire JDIA6_EBR,
	input wire JDIA7_EBR,
	input wire JDIA8_EBR,
	input wire JDIA9_EBR,
	input wire JDIB0_EBR,
	input wire JDIB10_EBR,
	input wire JDIB11_EBR,
	input wire JDIB12_EBR,
	input wire JDIB13_EBR,
	input wire JDIB14_EBR,
	input wire JDIB15_EBR,
	input wire JDIB16_EBR,
	input wire JDIB17_EBR,
	input wire JDIB1_EBR,
	input wire JDIB2_EBR,
	input wire JDIB3_EBR,
	input wire JDIB4_EBR,
	input wire JDIB5_EBR,
	input wire JDIB6_EBR,
	input wire JDIB7_EBR,
	input wire JDIB8_EBR,
	input wire JDIB9_EBR,

	input wire JOCEA_EBR,
	input wire JOCEB_EBR,
	input wire JRSTA_EBR,
	input wire JRSTB_EBR,
	input wire JWEA_EBR,
	input wire JWEB_EBR,

	output wire JDOB8_EBR,
	output wire JDOB16_EBR,
	output wire JDOB0_EBR,
	output wire JDOB9_EBR,
	output wire JDOB17_EBR,
	output wire JDOB1_EBR,
	output wire JDOB10_EBR,
	output wire JDOB2_EBR,
	output wire JDOB11_EBR,
	output wire JDOB3_EBR,
	output wire JDOB12_EBR,
	output wire JDOB4_EBR,
	output wire JDOB13_EBR,
	output wire JDOB5_EBR,
	output wire JDOB14_EBR,
	output wire JDOB6_EBR,
	output wire JDOB15_EBR,
	output wire JDOB7_EBR,
	output wire JDOA8_EBR,
	output wire JDOA16_EBR,
	output wire JDOA0_EBR,
	output wire JDOA9_EBR,
	output wire JDOA17_EBR,
	output wire JDOA1_EBR,
	output wire JDOA10_EBR,
	output wire JDOA2_EBR,
	output wire JDOA11_EBR,
	output wire JDOA3_EBR,
	output wire JDOA12_EBR,
	output wire JDOA4_EBR,
	output wire JDOA13_EBR,
	output wire JDOA5_EBR,
	output wire JDOA14_EBR,
	output wire JDOA6_EBR,
	output wire JDOA15_EBR,
	output wire JDOA7_EBR
);
	parameter INITVAL_00 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_01 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_02 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_03 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_04 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_05 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_06 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_07 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_08 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_09 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_0A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_0B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_0C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_0D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_0E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_0F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_10 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_11 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_12 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_13 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_14 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_15 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_16 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_17 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_20 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_21 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_22 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_23 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_24 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_25 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_26 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_27 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_28 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_29 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_2A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_2B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_2C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_2D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_2E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_2F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_30 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_31 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_32 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_33 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_34 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_35 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_36 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_37 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_38 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_39 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_3A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_3B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_3C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_3D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_3E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INITVAL_3F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_DATA = "STATIC";
	parameter CLKWMUX = "CLKW";
	parameter CLKRMUX = "CLKR";

	PDPW16KD PDPW16KD_inst (
		.BE({JADA12_EBR, JADA11_EBR, JADA10_EBR, JADA9_EBR}),
		.ADW({JADA13_EBR, JADA12_EBR, JADA11_EBR, JADA10_EBR, JADA9_EBR, JADA8_EBR, JADA7_EBR, JADA6_EBR, JADA5_EBR, JADA4_EBR, JADA3_EBR, JADA2_EBR, JADA1_EBR, JADA0_EBR}),
		.ADR({JADB13_EBR, JADB12_EBR, JADB11_EBR, JADB10_EBR, JADB9_EBR, JADB8_EBR, JADB7_EBR, JADB6_EBR, JADB5_EBR, JADB4_EBR, JADB3_EBR, JADB2_EBR, JADB1_EBR, JADB0_EBR}),
		.CSW({JCSA2_EBR, JCSA1_EBR, JCSA0_EBR}),
		.CSR({JCSB2_EBR, JCSB1_EBR, JCSB0_EBR}),
		.DI({JDIB17_EBR, JDIB16_EBR, JDIB15_EBR, JDIB14_EBR, JDIB13_EBR, JDIB12_EBR, JDIB11_EBR, JDIB10_EBR, JDIB9_EBR, JDIB8_EBR, JDIB7_EBR, JDIB6_EBR, JDIB5_EBR, JDIB4_EBR, JDIB3_EBR, JDIB2_EBR, JDIB1_EBR, JDIB0_EBR, JDIA17_EBR, JDIA16_EBR, JDIA15_EBR, JDIA14_EBR, JDIA13_EBR, JDIA12_EBR, JDIA11_EBR, JDIA10_EBR, JDIA9_EBR, JDIA8_EBR, JDIA7_EBR, JDIA6_EBR, JDIA5_EBR, JDIA4_EBR, JDIA3_EBR, JDIA2_EBR, JDIA1_EBR, JDIA0_EBR}),
		.DO({JDOB17_EBR, JDOB16_EBR, JDOB15_EBR, JDOB14_EBR, JDOB13_EBR, JDOB12_EBR, JDOB11_EBR, JDOB10_EBR, JDOB9_EBR, JDOB8_EBR, JDOB7_EBR, JDOB6_EBR, JDOB5_EBR, JDOB4_EBR, JDOB3_EBR, JDOB2_EBR, JDOB1_EBR, JDOB0_EBR, JDOA17_EBR, JDOA16_EBR, JDOA15_EBR, JDOA14_EBR, JDOA13_EBR, JDOA12_EBR, JDOA11_EBR, JDOA10_EBR, JDOA9_EBR, JDOA8_EBR, JDOA7_EBR, JDOA6_EBR, JDOA5_EBR, JDOA4_EBR, JDOA3_EBR, JDOA2_EBR, JDOA1_EBR, JDOA0_EBR}),
		.CLKW(JCLKA_EBR),
		.CLKR(JCLKB_EBR),
		.CEW(JCEA_EBR),
		.CER(JCEB_EBR),
		.OCER(JOCEB_EBR)
	);

endmodule

module PDPW16KD (
  input wire[13:0] ADR, // read address
  input wire[8:0] ADW, // write address
  input wire[3:0] BE, // ?
  input wire[2:0] CSW, // chip select write ?
  input wire[2:0] CSR, // chip select read ?
  output wire[35:0] DO, // dataout
  input wire CLKW, // write clock
  input wire[35:0] DI, // data in
  input wire CEW, // clock enable write
  input wire CLKR, // read clock
  input wire CER, //clock enable read
  input wire OCER // ?
);
  // 512 x 36 memory;

  reg[35:0] memory[511:0];
  reg[35:0] next_memory[511:0];

  reg[35:0] next_DO, DO_reg;

  integer i, i2;

  always @ (*) begin
    for (i = 0; i < 512; i = i + 1) begin
      next_memory[i] = memory[i];
    end
    if (CEW && BE[0]) begin
      next_memory[ADW] = DI;
    end
  end

  always @ (posedge CLKW) begin
    for (i2 = 0; i2 < 512; i2 = i2 + 1) begin
      memory[i2] <= next_memory[i2];
    end
  end

  always @ (*) begin
    next_DO = 36'b0;
    if (CER) begin
      next_DO = memory[ADR[13:5]];
    end
  end

  always @ (posedge CLKR) begin
    DO_reg <= next_DO;
  end

  assign DO = DO_reg;

endmodule